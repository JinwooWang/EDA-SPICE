
V1 1 0 sin(0 1 1)
R1 1 2 0.01
D1 2 0 D1N4148
.TRAN 1ns 5ns
