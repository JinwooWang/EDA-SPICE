
M2 2 1 0 2 MOD1 W=2 L=1
V1 1 0 1.5
V2 2 0 1.5
.MODEL MOD1 NMOS
.MODEL MOD2 PMOS
.DC V2 0 5 0.1
