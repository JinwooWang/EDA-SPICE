*elmore
v1 1 0 pulse(0 3 2ns 2ns 2ns 15ns 30ns)
R1 1 2 1
C1 2 0 2
R2 2 3 1
C2 3 0 2
R3 2 4 1
C3 4 0 2
R4 4 5 1
C4 5 0 2
R5 4 6 1
C6 6 0 2

.tran 1ns 35ns
.end
