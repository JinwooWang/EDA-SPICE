
Vs 1 0 5
R1 1 2 5
L1 1 2 4
C1 2 0 5
.TRAN 1NS 30NS
