opamp
Vdd 1 0 1.8
R1 1 2 50k
M1 2 2 0 0 MOD1 W=1 L=1
M2 4 4 1 1 MOD2 W=4 L=1
M3 5 4 1 1 MOD2 W=4 L=1
M4 4 8 3 3 MOD1 W=10 L=1
M5 5 9 3 3 MOD1 W=10 L=1
M6 3 2 0 0 MOD1 W=1 L=1
M7 7 5 1 1 MOD2 W=4 L=1
M8 7 2 0 0 MOD1 W=6 L=1
Cc 5 6 200f
R2 6 7 10K
Vm 8 0 1.8
Vp 9 0 sin(0 1 1)
Cp 7 0 10p
.TRAN 1ns 5ns
.MODEL MOD1 NMOS
.MODEL MOD2 PMOS

.END
